module shurf

struct StaticFile {
	path string
	size usize
}
