module shurf

pub type Handler = fn (ctx Context) ?
