module shurf

pub type Handler<U> = fn (ctx Context<U>) ?
