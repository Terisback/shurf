module shurf

pub struct Config {
pub mut:
	app_name string
}
