module shurf

struct Pool {
}
