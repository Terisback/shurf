module pevo
