module shurf
