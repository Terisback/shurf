module utils

[noinit]
pub struct ErrOutOfBounds {
pub:
	msg  string = 'out of bounds'
	code int    = 1
}
